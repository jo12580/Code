** Profile: "SCHEMATIC2-2"  [ G:\030\12.7\13_4-PSpiceFiles\SCHEMATIC2\2.sim ] 

** Creating circuit file "2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10U 0 
.OPTIONS ADVCONV
.OPTIONS DIGINITSTATE= 0
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC2.net" 


.END
