** Profile: "Voltage as scanning variable-2-DC-R2"  [ D:\Software\Capture_PSpice\Project\DC scan analysis\DC scan analysis-PSpiceFiles\Voltage as scanning variable\2-DC-R2.sim ] 

** Creating circuit file "2-DC-R2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN PARAM rvar 1k 10k 10 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Voltage as scanning variable.net" 


.END
