** Profile: "��̬���������-007"  [ D:\Software\Capture_PSpice\Project\Static operating point analysis circuit\Static operating point analysis circuit-PSpiceFiles\��̬���������\007.sim ] 

** Creating circuit file "007.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.OP
.OPTIONS ADVCONV
.OPTIONS ITL2= 200
.OPTIONS ITL4= 100
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\��̬���������.net" 


.END
