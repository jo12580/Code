** Profile: "SCHEMATIC2-2"  [ D:\Software\Capture_PSpice\Project\PSPICE06\06-PSpiceFiles\SCHEMATIC2\2.sim ] 

** Creating circuit file "2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../06-pspicefiles/06.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10m 0 0.01m 
.FOUR 1k 9 V([OUT]) 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC2.net" 


.END
