** Profile: "schematic2-page2_tran"  [ D:\Software\Capture_PSpice\Project\Electronic circuit design\exam_1-pspicefiles\schematic2\page2_tran.sim ] 

** Creating circuit file "page2_tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 15m 0 0.01m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\schematic2.net" 


.END
