** Profile: "Digital_analog_mixing-4"  [ D:\Software\Capture_PSpice\Project\Digital analog hybrid circuit\Digital signal source-PSpiceFiles\Digital_analog_mixing\4.sim ] 

** Creating circuit file "4.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 50u 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Digital_analog_mixing.net" 


.END
