** Profile: "Exponential_signal_source-4"  [ D:\Software\Capture_PSpice\Project\Transient analysis and Fourier analysis\Transient analysis and Fourier analysis-PSpiceFiles\Exponential_signal_source\4.sim ] 

** Creating circuit file "4.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 20ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Exponential_signal_source.net" 


.END
