** Profile: "SCHEMATIC1-3"  [ D:\Software\Capture_PSpice\Project\Transmission scan analysis\Transmission scan analysis-PSpiceFiles\SCHEMATIC1\3.sim ] 

** Creating circuit file "3.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_VCC2 0 10 0.01 
.STEP LIN I_IBB2 0 100u 10u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
