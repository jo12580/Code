** Profile: "SCHEMATIC1-3"  [ G:\030\11.23\23-pspicefiles\schematic1\3.sim ] 

** Creating circuit file "3.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ad627a/ad627a.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "G:\030\11.23\AD627A\AD627A.lib" 
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 1 0.1 100k
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
