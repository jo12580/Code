** Profile: "Transient_analysis-Transient_analysis"  [ D:\Software\Capture_PSpice\Project\Transient analysis and Fourier analysis\Transient analysis and Fourier analysis-PSpiceFiles\Transient_analysis\Transient_analysis.sim ] 

** Creating circuit file "Transient_analysis.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10u 0 0.001 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Transient_analysis.net" 


.END
